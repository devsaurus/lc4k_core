
library ieee;
use ieee.std_logic_1164.all;

entity reg_pipe_cpld is

  port (
    i_clk : in  std_logic;
    i_ce  : in  std_logic;
    i_res : in  std_logic;
    i_d   : in  std_logic_vector(7 downto 0);
    o_d   : out std_logic_vector(7 downto 0);
    o_or  : out std_logic
  );

end;

architecture struct of reg_pipe_cpld is

  constant c_fusemap : std_logic_vector(0 to 17200-1) :=
"1111100011000110001100011111110001111111000111111100010000111111111111111111111111111111110000110001100011000110001000011111110001111111000111111111111000111111111111111111" &
"1101100011000110001100011111110001111111000111111100011000111111111111111111111111111111000000110001100011000110001100011111110001111111000111111111111000111111111111111111" &
"1111100011000100001100011111110001111111000111111100011000111111111111111111111111111111110000110001100010000110001100011111110001111111000111111111111000111111111111111111" &
"1101100011000110001100011111110001111111000111111100011000111111111111111111111111111111000000110001100011000110001100011111110001111111000111111111111000111111111111111111" &
"1101100011000110001100011111110001111111000111111000011000111111111111111111111111111111010000110001100011000110001100011111110001111110000111111111111000111111111111111111" &
"1111100011000110001100011111110001111111000111111100011000111111111111111111111111111111100000110001100011000110001100011111110001111111000111111111111000111111111111111111" &
"1101100011000110001100011111110001111110000111111100011000111111111111111111111111111101110000110001100011000110001100011111010001111111000111111111111000111111111111111111" &
"1111100011000110001100011111110001111111000111111100011000111111111111111111111111111111110000110001100011000110001100011111110001111111000111111111111000111111111111111111" &
"1111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111" &
"1101111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1101111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1101111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111101111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1010111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111011111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111011" &
"1011111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1101111111111111111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111011110111101111011111111101111111110111111111011110111111111111111111111111111111111111111011110111101111011110111111111011111111101111111111111101111111111111111111111" &
"1010111101111011110111111111011111111101111111110111101111111111111111111111111111111110111111101111011110111101111011111111101111111110111111111111110111111111111111111111" &
"1111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1101111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1101111111111111111111111111011111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111111111011111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1101111111111111110111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111110111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111101111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111110111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111101111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111101111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111111011111111101111111110111111110111111111111111111111111111111111111011111111001111111100111111111011111111101111111111111111110111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111111011111111101111111110111111110111111111111111111111111111111111111011111111001111111100111111111011111111101111111111111111110111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111111011111111101111111110111111110111111111111111111111111111111111111011111111001111111100111111111011111111101111111111111111110111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111101111111100111111111011111111001111111100111111111111110111111111011111111101111111110111111111011111111100111111111011111111001111111" &
"1111111001111111100111111111011111111101111111101111111110011111111001111111100111111111111110011111111011111111110111111110011111111001111111100111111110011111111001111111" &
"1111111001111111100111111111011111111001111111100111111110011111111001111111100111111111111110111111111101111111100111111110011111111001111111100111111110011111111001111111" &
"1111111001111111100111111110011111111001111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111011" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111111111111111111111111111111111111111111111111110111111111111111111110111111110011111111001111111100111111110011111111011111111"
;

  signal ncon : std_logic;
  signal pu, pd, kp : std_logic;

  signal d_out  : std_logic_vector(o_d'range);
  signal or_out : std_logic;

begin

  cpld_b : entity work.lc4032x_tqfp48_core
    generic map (
      g_fusemap => c_fusemap
    )
    port map (
      i_2    => i_ce,
      o_2    => open,
      oe_2   => open,
      i_3    => i_res,
      o_3    => open,
      oe_3   => open,
      i_4    => i_d(0),
      o_4    => open,
      oe_4   => open,
      i_7    => i_d(1),
      o_7    => open,
      oe_7   => open,
      i_8    => i_d(2),
      o_8    => open,
      oe_8   => open,
      i_9    => i_d(3),
      o_9    => open,
      oe_9   => open,
      i_10   => i_d(4),
      o_10   => open,
      oe_10  => open,
      i_14   => i_d(5),
      o_14   => open,
      oe_14  => open,
      i_15   => i_d(6),
      o_15   => open,
      oe_15  => open,
      i_16   => i_d(7),
      o_16   => open,
      oe_16  => open,
      i_17   => ncon,
      o_17   => open,
      oe_17  => open,
      i_18   => i_clk,
      i_19   => ncon,
      i_20   => d_out(0),
      o_20   => d_out(0),
      oe_20  => open,
      i_21   => d_out(1),
      o_21   => d_out(1),
      oe_21  => open,
      i_22   => d_out(2),
      o_22   => d_out(2),
      oe_22  => open,
      i_23   => d_out(3),
      o_23   => d_out(3),
      oe_23  => open,
      i_24   => d_out(4),
      o_24   => d_out(4),
      oe_24  => open,
      i_26   => d_out(5),
      o_26   => d_out(5),
      oe_26  => open,
      i_27   => d_out(6),
      o_27   => d_out(6),
      oe_27  => open,
      i_28   => d_out(7),
      o_28   => d_out(7),
      oe_28  => open,
      i_31   => ncon,
      o_31   => open,
      oe_31  => open,
      i_32   => ncon,
      o_32   => open,
      oe_32  => open,
      i_33   => ncon,
      o_33   => open,
      oe_33  => open,
      i_34   => ncon,
      o_34   => open,
      oe_34  => open,
      i_38   => ncon,
      o_38   => open,
      oe_38  => open,
      i_39   => ncon,
      o_39   => open,
      oe_39  => open,
      i_40   => ncon,
      o_40   => open,
      oe_40  => open,
      i_41   => ncon,
      o_41   => open,
      oe_41  => open,
      i_42   => ncon,
      i_43   => ncon,
      i_44   => or_out,
      o_44   => or_out,
      oe_44  => open,
      i_45   => ncon,
      o_45   => open,
      oe_45  => open,
      i_46   => ncon,
      o_46   => open,
      oe_46  => open,
      i_47   => ncon,
      o_47   => open,
      oe_47  => open,
      i_48   => ncon,
      o_48   => open,
      oe_48  => open,
      --
      o_pu => pu,
      o_pd => pd,
      o_kp => kp
    );

  ncon <= '1' when pu = '1' else
          '0' when pd = '1' else
          '1';

  o_d  <= d_out;
  o_or <= or_out;

end;
