
library ieee;
use ieee.std_logic_1164.all;

entity xor_in_cpld is

  port (
    i_xor : in  std_logic_vector(29 downto 0);
    o_out : out std_logic
  );

end;

architecture struct of xor_in_cpld is

  constant c_fusemap : std_logic_vector(0 to 17200-1) :=
"1111111111111111111111111111111111111111111111111111011111111111000011111111111111101111111111111111111111111111111111111111111111111111000111111111111000111111111111111011" &
"1101111111111111111111111111111111111111111111111111011111111110100011111111111111101111111111111111111111111111111111111111111111111111000111111111111000111111111111111011" &
"1111111111100111111111111111111111111111111111111111011111111111100011111111111111101111111111111111111111111111111111111111111111111110000111111111111000111111111111111011" &
"1011111110011111111111111111111111111111111111111111011111111111100011111111111111101111011111111111111111111111111111111111111111111101000111111111111000111111111111111011" &
"1111111111111111111111111111111111111111111111111010011111111111100011111111111111101111111111111001111111111111111111111111111111111111000111111111111000111111111111111011" &
"0111111111111111111111111111111111111111111111110101011111111111100011111111111111101111011111100111111111111111111111111111111111111111000111111111111000111111111111111011" &
"1111111111111111111111111111111111111111111111111111011111111111100011111111111111101111011111110101111111111111111111111111111111111111000111111111111000111111111111111011" &
"1011111111111111111111111111011111111111111111111111011111111111100011111111111111101111111111101011111111111111111111111111111111111111000111111111111000111111111111111011" &
"1101111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111" &
"1111111111111111111111111111111111111111111111110011111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111101111111111111111111111" &
"1101111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111011111111111111111111101111111111111111111111111111111111111011111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111010111111111111111111111111111111111111111111101111111111111111111111111111101011111111111111111111111111111111111111111111111111111" &
"0111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111100111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111" &
"0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111" &
"1111111111111111110111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111101011111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111100111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"0111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111111111111111111111111110011111111111111111111111111111111111111111111111111111101111111111111111111111111111110011111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111" &
"1011111111111111111111111111111001111111111111111111111111111111111111111111111111111101111111111111111111111111111100111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111" &
"1011111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111001111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101101111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111001111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111101111111111111111111111" &
"0111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111100111111111111111111111111111111111111111111111" &
"0111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"0111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"0111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111101101111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"0111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111010111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1011111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111101111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111010111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111001111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111" &
"0111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111101111111110111111111011111111101111111111111111111111111111111111111111111111111111111011111111101111111110111111111011111111111111111111111111111111111111111111111" &
"1111111101111111110111111111011111111101111111110111111111111111111011111111111111111111111111011111111101111111110111111111011111111101111111111111111110111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111101111111110111111111011111111101111111110111111111111111111011111111111111111111111111011111111101111111110111111111011111111101111111111111111110111111111111111111" &
"1111111101111111110111111111011111111101111111110111111111111111111011111111111111111111111111011111111101111111110111111111011111111101111111111111111110111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111011111111101111111110111111111011111111101111111110011111111101111111100111111111111111111111111011111111101111111110111111111011111111100111111111011111111001111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111101111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111"
;

  signal ncon : std_logic;
  signal pu, pd, kp : std_logic;

  signal out_s : std_logic;

begin

  cpld_b : entity work.lc4032x_tqfp48_core
    generic map (
      g_fusemap => c_fusemap
    )
    port map (
      i_2    => i_xor(0),
      o_2    => open,
      oe_2   => open,
      i_3    => i_xor(1),
      o_3    => open,
      oe_3   => open,
      i_4    => i_xor(2),
      o_4    => open,
      oe_4   => open,
      i_7    => i_xor(3),
      o_7    => open,
      oe_7   => open,
      i_8    => i_xor(4),
      o_8    => open,
      oe_8   => open,
      i_9    => i_xor(5),
      o_9    => open,
      oe_9   => open,
      i_10   => i_xor(6),
      o_10   => open,
      oe_10  => open,
      i_14   => i_xor(7),
      o_14   => open,
      oe_14  => open,
      i_15   => i_xor(8),
      o_15   => open,
      oe_15  => open,
      i_16   => i_xor(9),
      o_16   => open,
      oe_16  => open,
      i_17   => i_xor(10),
      o_17   => open,
      oe_17  => open,
      i_18   => ncon,
      i_19   => ncon,
      i_20   => i_xor(11),
      o_20   => open,
      oe_20  => open,
      i_21   => i_xor(12),
      o_21   => open,
      oe_21  => open,
      i_22   => i_xor(13),
      o_22   => open,
      oe_22  => open,
      i_23   => i_xor(14),
      o_23   => open,
      oe_23  => open,
      i_24   => i_xor(15),
      o_24   => open,
      oe_24  => open,
      i_26   => i_xor(16),
      o_26   => open,
      oe_26  => open,
      i_27   => i_xor(17),
      o_27   => open,
      oe_27  => open,
      i_28   => i_xor(18),
      o_28   => open,
      oe_28  => open,
      i_31   => i_xor(19),
      o_31   => open,
      oe_31  => open,
      i_32   => i_xor(20),
      o_32   => open,
      oe_32  => open,
      i_33   => i_xor(21),
      o_33   => open,
      oe_33  => open,
      i_34   => i_xor(22),
      o_34   => open,
      oe_34  => open,
      i_38   => i_xor(23),
      o_38   => open,
      oe_38  => open,
      i_39   => i_xor(24),
      o_39   => open,
      oe_39  => open,
      i_40   => i_xor(25),
      o_40   => open,
      oe_40  => open,
      i_41   => ncon,
      o_41   => open,
      oe_41  => open,
      i_42   => ncon,
      i_43   => ncon,
      i_44   => out_s,
      o_44   => out_s,
      oe_44  => open,
      i_45   => i_xor(26),
      o_45   => open,
      oe_45  => open,
      i_46   => i_xor(27),
      o_46   => open,
      oe_46  => open,
      i_47   => i_xor(28),
      o_47   => open,
      oe_47  => open,
      i_48   => i_xor(29),
      o_48   => open,
      oe_48  => open,
      --
      o_pu => pu,
      o_pd => pd,
      o_kp => kp
    );

  ncon <= '1' when pu = '1' else
          '0' when pd = '1' else
          '1';

  o_out <= out_s;

end;
