
library ieee;
use ieee.std_logic_1164.all;

entity bclk_set_res_cpld is

  port (
    i_clk_a    : in  std_logic;
    i_clk_b    : in  std_logic;
    i_setres_a : in  std_logic;
    i_setres_b : in  std_logic;
    i_setres_c : in  std_logic;
    i_setres_d : in  std_logic;
    i_din      : in  std_logic_vector(3 downto 0);
    o_dout     : out std_logic_vector(3 downto 0)
  );

end;

architecture struct of bclk_set_res_cpld is

  constant c_fusemap : std_logic_vector(0 to 17200-1) :=
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111101001111110100111111010011111100001111111111111111111111111101001111111111011" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111110100111111010011111100001111111111111111111111111101001111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111101111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111011111111111111111111111111111111111111111111111110111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111011" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111011111111111111111111111111111111111111111111111110111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111110111111111011111111111111111111111111111011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111110111111111111111111111111111111111111111011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111110111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111011111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111110111111111111111111111111111111111111111011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111011111111101111111110111111111111111111111111111111111111111011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111011111111101111111110111111111001111111100111111110011111111101111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111101111111" &
"1111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111110011111111001111111100111111110011111111001111111100111111110011111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111011111111001111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111011111111001111001" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111011111111001111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111110111111110011111111001111111100111111110011111111001111111"
;

  signal ncon : std_logic;
  signal pu, pd, kp : std_logic;

  signal dout : std_logic_vector(o_dout'range);

begin

  cpld_b : entity work.lc4032zc_tqfp48_core
    generic map (
      g_fusemap => c_fusemap
    )
    port map (
      i_2    => i_din(0),
      o_2    => open,
      oe_2   => open,
      i_3    => i_din(1),
      o_3    => open,
      oe_3   => open,
      i_4    => i_din(2),
      o_4    => open,
      oe_4   => open,
      i_7    => i_din(3),
      o_7    => open,
      oe_7   => open,
      i_8    => i_setres_a,
      o_8    => open,
      oe_8   => open,
      i_9    => i_setres_b,
      o_9    => open,
      oe_9   => open,
      i_10   => i_setres_c,
      o_10   => open,
      oe_10  => open,
      i_14   => i_setres_d,
      o_14   => open,
      oe_14  => open,
      i_15   => dout(0),
      o_15   => dout(0),
      oe_15  => open,
      i_16   => dout(1),
      o_16   => dout(1),
      oe_16  => open,
      i_17   => dout(2),
      o_17   => dout(2),
      oe_17  => open,
      i_18   => i_clk_a,
      i_19   => i_clk_b,
      i_20   => ncon,
      o_20   => open,
      oe_20  => open,
      i_21   => ncon,
      o_21   => open,
      oe_21  => open,
      i_22   => ncon,
      o_22   => open,
      oe_22  => open,
      i_23   => ncon,
      o_23   => open,
      oe_23  => open,
      i_24   => ncon,
      o_24   => open,
      oe_24  => open,
      i_26   => ncon,
      o_26   => open,
      oe_26  => open,
      i_27   => ncon,
      o_27   => open,
      oe_27  => open,
      i_28   => ncon,
      o_28   => open,
      oe_28  => open,
      i_31   => ncon,
      o_31   => open,
      oe_31  => open,
      i_32   => ncon,
      o_32   => open,
      oe_32  => open,
      i_33   => ncon,
      o_33   => open,
      oe_33  => open,
      i_34   => ncon,
      o_34   => open,
      oe_34  => open,
      i_38   => ncon,
      o_38   => open,
      oe_38  => open,
      i_39   => ncon,
      o_39   => open,
      oe_39  => open,
      i_40   => ncon,
      o_40   => open,
      oe_40  => open,
      i_41   => ncon,
      o_41   => open,
      oe_41  => open,
      i_42   => ncon,
      i_43   => ncon,
      i_44   => ncon,
      o_44   => open,
      oe_44  => open,
      i_45   => dout(3),
      o_45   => dout(3),
      oe_45  => open,
      i_46   => ncon,
      o_46   => open,
      oe_46  => open,
      i_47   => ncon,
      o_47   => open,
      oe_47  => open,
      i_48   => ncon,
      o_48   => open,
      oe_48  => open,
      --
      o_pu => pu,
      o_pd => pd,
      o_kp => kp
    );

  ncon <= '1' when pu = '1' else
          '0' when pd = '1' else
          '1';

  o_dout <= dout;

end;
