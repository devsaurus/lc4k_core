
library ieee;
use ieee.std_logic_1164.all;

entity oe_cpld is

  port (
    i_clk : in  std_logic;
    i_res : in  std_logic;
    i_oe  : in  std_logic;
    i_d   : in  std_logic_vector(7 downto 0);
    o_d   : out std_logic_vector(7 downto 0)
  );

end;

architecture struct of oe_cpld is

  constant c_fusemap : std_logic_vector(0 to 35600-1) :=
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111000011111100001111110001111110000011111111111111110000111111111111111111111111101111111111111000011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100001111110001111111000011111111111111110000111111111111111111111111111111111111111100011111111111100001111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111101111111110111111111111111111101111111111111111111111111111111111111111111111101111111111011111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111101111111110111111111111111111101111111111111111111111111111111111111111111111101111111111011111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111110011111111001111111100111111110011111111001111111100111111110011111111001111110111111111100111111110011111111001111111100111111110011111111001111111100111111110011111111111111111001111111100111111110011111111001111111100111111110011111111001111111100111111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111101111111110111111111111111111101111111111111111111111111111111111111111111111101111111111011111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110" &
"11111111110011111111001111111100111111110011111111001111111100111111110011111111001111111111111111100111111111111111111111111111101111111111011111111001111111100111111110011111111111111111001111111110111111111111111111001111111100111111111011111111001111111100111111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"11111111110011111111001111111100111111110011111111001111111100111111110011111111001111111111111111101111111110011111111001111111100111111111011111111011111111100111111110011111111111111111101111111100111111110011111111001111111100111111110011111111001111111100111111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"11111111110011111111001111111100111111110011111111001111111100111111110011111111001111111111111111101111111110011111111001111111100111111110011111111011111111100111111110011111111111111111001111111100111111110111111111001111111100111111110011111111001111111100111111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111011111111111111111110111111111101111111111111111111111111111111111111011111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111011111111111111111110111111111101111111111111111111111111111111111111011111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111111111111111111111110111111111101111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111011111111111111111110111111111101111111111111111111111111111111111111011111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111" &
"11111111011111111111011011111101101111110011111101111011110111101111011110111101111011111111111110110111111110111111111011011110111111111110111111101101111110111111111111111111111111111111011111110111101111110011111101111111110111101111011110111101111011110111101111111111111110011111111011111111101111111110111111111011111110111101111011111111111111111111"
  ;

  signal ncon : std_logic;

  signal d_out, d_oe : std_logic_vector(o_d'range);

begin

  cpld_b : entity work.lc4064ze_csbga64_core
    generic map (
      g_fusemap => c_fusemap
    )
    port map (
      i_A1   => i_res,
      o_A1   => open,
      oe_A1  => open,
      pu_A1  => open,
      pd_A1  => open,
      kp_A1  => open,
      i_A2   => i_d(0),
      o_A2   => open,
      oe_A2  => open,
      pu_A2  => open,
      pd_A2  => open,
      kp_A2  => open,
      i_A3   => i_d(1),
      o_A3   => open,
      oe_A3  => open,
      pu_A3  => open,
      pd_A3  => open,
      kp_A3  => open,
      i_A4   => i_clk,
      pu_A4  => open,
      pd_A4  => open,
      kp_A4  => open,
      i_A5   => i_d(2),
      o_A5   => open,
      oe_A5  => open,
      pu_A5  => open,
      pd_A5  => open,
      kp_A5  => open,
      i_A6   => i_d(3),
      o_A6   => open,
      oe_A6  => open,
      pu_A6  => open,
      pd_A6  => open,
      kp_A6  => open,
      i_A7   => i_d(4),
      o_A7   => open,
      oe_A7  => open,
      pu_A7  => open,
      pd_A7  => open,
      kp_A7  => open,
      i_A8   => i_d(5),
      o_A8   => open,
      oe_A8  => open,
      pu_A8  => open,
      pd_A8  => open,
      kp_A8  => open,
      i_B1   => i_d(6),
      o_B1   => open,
      oe_B1  => open,
      pu_B1  => open,
      pd_B1  => open,
      kp_B1  => open,
      i_B3   => i_d(7),
      o_B3   => open,
      oe_B3  => open,
      pu_B3  => open,
      pd_B3  => open,
      kp_B3  => open,
      i_B4   => i_oe,
      o_B4   => open,
      oe_B4  => open,
      pu_B4  => open,
      pd_B4  => open,
      kp_B4  => open,
      i_B5   => ncon,
      o_B5   => open,
      oe_B5  => open,
      pu_B5  => open,
      pd_B5  => open,
      kp_B5  => open,
      i_B6   => ncon,
      o_B6   => open,
      oe_B6  => open,
      pu_B6  => open,
      pd_B6  => open,
      kp_B6  => open,
      i_B7   => ncon,
      o_B7   => open,
      oe_B7  => open,
      pu_B7  => open,
      pd_B7  => open,
      kp_B7  => open,
      i_C1   => ncon,
      o_C1   => open,
      oe_C1  => open,
      pu_C1  => open,
      pd_C1  => open,
      kp_C1  => open,
      i_C2   => ncon,
      o_C2   => open,
      oe_C2  => open,
      pu_C2  => open,
      pd_C2  => open,
      kp_C2  => open,
      i_C3   => ncon,
      o_C3   => open,
      oe_C3  => open,
      pu_C3  => open,
      pd_C3  => open,
      kp_C3  => open,
      i_C4   => ncon,
      pu_C4  => open,
      pd_C4  => open,
      kp_C4  => open,
      i_C5   => ncon,
      o_C5   => open,
      oe_C5  => open,
      pu_C5  => open,
      pd_C5  => open,
      kp_C5  => open,
      i_C7   => ncon,
      o_C7   => open,
      oe_C7  => open,
      pu_C7  => open,
      pd_C7  => open,
      kp_C7  => open,
      i_C8   => ncon,
      o_C8   => open,
      oe_C8  => open,
      pu_C8  => open,
      pd_C8  => open,
      kp_C8  => open,
      i_D1   => ncon,
      o_D1   => open,
      oe_D1  => open,
      pu_D1  => open,
      pd_D1  => open,
      kp_D1  => open,
      i_D2   => ncon,
      o_D2   => open,
      oe_D2  => open,
      pu_D2  => open,
      pd_D2  => open,
      kp_D2  => open,
      i_D3   => ncon,
      o_D3   => open,
      oe_D3  => open,
      pu_D3  => open,
      pd_D3  => open,
      kp_D3  => open,
      i_D7   => ncon,
      o_D7   => open,
      oe_D7  => open,
      pu_D7  => open,
      pd_D7  => open,
      kp_D7  => open,
      i_D8   => ncon,
      o_D8   => open,
      oe_D8  => open,
      pu_D8  => open,
      pd_D8  => open,
      kp_D8  => open,
      i_E1   => ncon,
      o_E1   => open,
      oe_E1  => open,
      pu_E1  => open,
      pd_E1  => open,
      kp_E1  => open,
      i_E2   => ncon,
      o_E2   => open,
      oe_E2  => open,
      pu_E2  => open,
      pd_E2  => open,
      kp_E2  => open,
      i_E6   => ncon,
      o_E6   => open,
      oe_E6  => open,
      pu_E6  => open,
      pd_E6  => open,
      kp_E6  => open,
      i_E7   => ncon,
      o_E7   => open,
      oe_E7  => open,
      pu_E7  => open,
      pd_E7  => open,
      kp_E7  => open,
      i_E8   => ncon,
      o_E8   => open,
      oe_E8  => open,
      pu_E8  => open,
      pd_E8  => open,
      kp_E8  => open,
      i_F1   => ncon,
      o_F1   => open,
      oe_F1  => open,
      pu_F1  => open,
      pd_F1  => open,
      kp_F1  => open,
      i_F2   => ncon,
      o_F2   => open,
      oe_F2  => open,
      pu_F2  => open,
      pd_F2  => open,
      kp_F2  => open,
      i_F3   => ncon,
      o_F3   => open,
      oe_F3  => open,
      pu_F3  => open,
      pd_F3  => open,
      kp_F3  => open,
      i_F5   => ncon,
      o_F5   => open,
      oe_F5  => open,
      pu_F5  => open,
      pd_F5  => open,
      kp_F5  => open,
      i_F6   => ncon,
      o_F6   => open,
      oe_F6  => open,
      pu_F6  => open,
      pd_F6  => open,
      kp_F6  => open,
      i_F7   => ncon,
      o_F7   => open,
      oe_F7  => open,
      pu_F7  => open,
      pd_F7  => open,
      kp_F7  => open,
      i_F8   => ncon,
      o_F8   => open,
      oe_F8  => open,
      pu_F8  => open,
      pd_F8  => open,
      kp_F8  => open,
      i_G1   => ncon,
      o_G1   => open,
      oe_G1  => open,
      pu_G1  => open,
      pd_G1  => open,
      kp_G1  => open,
      i_G2   => ncon,
      o_G2   => open,
      oe_G2  => open,
      pu_G2  => open,
      pd_G2  => open,
      kp_G2  => open,
      i_G3   => ncon,
      o_G3   => open,
      oe_G3  => open,
      pu_G3  => open,
      pd_G3  => open,
      kp_G3  => open,
      i_G4   => ncon,
      pu_G4  => open,
      pd_G4  => open,
      kp_G4  => open,
      i_G5   => d_out(0),
      o_G5   => d_out(0),
      oe_G5  => d_oe(0),
      pu_G5  => open,
      pd_G5  => open,
      kp_G5  => open,
      i_G6   => d_out(1),
      o_G6   => d_out(1),
      oe_G6  => d_oe(1),
      pu_G6  => open,
      pd_G6  => open,
      kp_G6  => open,
      i_G7   => d_out(2),
      o_G7   => d_out(2),
      oe_G7  => d_oe(2),
      pu_G7  => open,
      pd_G7  => open,
      kp_G7  => open,
      i_G8   => d_out(3),
      o_G8   => d_out(3),
      oe_G8  => d_oe(3),
      pu_G8  => open,
      pd_G8  => open,
      kp_G8  => open,
      i_H2   => d_out(4),
      o_H2   => d_out(4),
      oe_H2  => d_oe(4),
      pu_H2  => open,
      pd_H2  => open,
      kp_H2  => open,
      i_H3   => d_out(5),
      o_H3   => d_out(5),
      oe_H3  => d_oe(5),
      pu_H3  => open,
      pd_H3  => open,
      kp_H3  => open,
      i_H4   => d_out(6),
      o_H4   => d_out(6),
      oe_H4  => d_oe(6),
      pu_H4  => open,
      pd_H4  => open,
      kp_H4  => open,
      i_H5   => ncon,
      pu_H5  => open,
      pd_H5  => open,
      kp_H5  => open,
      i_H6   => d_out(7),
      o_H6   => d_out(7),
      oe_H6  => d_oe(7),
      pu_H6  => open,
      pd_H6  => open,
      kp_H6  => open,
      i_H7   => ncon,
      o_H7   => open,
      oe_H7  => open,
      pu_H7  => open,
      pd_H7  => open,
      kp_H7  => open,
      --
      i_oscclk => '0'
    );

  ncon <= '1';

  oe_gen: for idx in o_d'range generate
    o_d(idx) <= d_out(idx) when d_oe(idx) = '1' else 'Z';
  end generate;

end;
